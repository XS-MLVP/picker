module {{__TOP_MODULE_NAME__}}_top;

{{__LOGIC_PIN_DECLARATION__}}

  {{__SOURCE_MOUDLE_NAME__}} {{__TOP_MODULE_NAME__}} (
{{__PIN_CONNECT__}}
  );

{{__DPI_FUNCTION_EXPORT__}}

{{__DPI_FUNCTION_IMPLEMENT__}}

{{__SV_DUMP_WAVE__}}

endmodule
