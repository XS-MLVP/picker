module {{__TOP_MODULE_NAME__}}_top;

{{__WIRE_PIN_DECLARATION__}}

{{__SOURCE_MODULE_NAME__}} {{__TOP_MODULE_NAME__}} (
{{__PIN_CONNECT__}}
  );
endmodule
