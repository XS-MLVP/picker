module {{__TOP_MODULE_NAME__}}_top(
    {{__INOUT_PIN_DECLARATION__}}
);

{{__LOGIC_PIN_DECLARATION__}}

{{__INOUT_PIN_ASSIGNMENT__}}

{{__INNER_MODULES__}}

{{__DPI_FUNCTION_EXPORT__}}

{{__DPI_FUNCTION_IMPLEMENT__}}

{{__SV_DUMP_WAVE__}}

{{__EXTEND_SV__}}

endmodule
