module {{__TOP_MODULE_NAME__}}_top;

{{__WIRE_PIN_DECLARATION__}}

{{__INNER_MODULES__}}

endmodule
