module Testmodule (
    input clk,
    input rst,
    input [31:0] addr,
    input [31:0] data_in,
    output [31:0] data_out,
    input [3:0]  cmd
);

endmodule;